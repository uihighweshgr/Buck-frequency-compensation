C:\USERS\USER\DOWNLOADS\BUCK_COMPENSATE_TYPEIII_CLOSELOOP.CIR/CONFIG 1/SETUP1
*#SAVE V(1) V(5) V(6) @VI[I] @VI[P] V(11) V(7) V(4)
*#SAVE V(3) @VREF[I] @VREF[P] V(2) V(8) @VIO[I] @VIO[P] V(14)
*#SAVE V(9)
*#ALIAS VO  V(3)
*#VIEW  AC VO
*#VIEW  AC PH_VO = PHASE(VO)
*#VIEW  TRAN VO
*#ALIAS VD  V(11)
*#VIEW  AC VD
*#VIEW  AC PH_VD = PHASE(VD)
*#VIEW  TRAN VD
*#ALIAS VIO  V(6)
*#VIEW  AC VIO
*#VIEW  AC PH_VIO = PHASE(VIO)
*#VIEW  TRAN VIO
*#ALIAS VGVG  V(5)
*#VIEW  AC VGVG
*#VIEW  AC PH_VGVG = PHASE(VGVG)
*#VIEW  TRAN VGVG
*#ALIAS VGVD  V(7)
*#VIEW  AC VGVD
*#VIEW  AC PH_VGVD = PHASE(VGVD)
*#VIEW  TRAN VGVD
*#ALIAS VIO2  V(4)
*#VIEW  AC VIO2
*#VIEW  AC PH_VIO2 = PHASE(VIO2)
*#VIEW  TRAN VIO2
*#ALIAS VI  V(1)
*#VIEW  AC VI
*#VIEW  AC PH_VI = PHASE(VI)
*#VIEW  TRAN VI
.AC DEC 10 1 1G
.TRAN 1N 16M
.OPTIONS ABSTOL=10N ITL4=200
.OPTIONS RELTOL=0.01 VNTOL=10U
.OPTIONS ACCT
.OPTIONS BYPASS=0
.PRINT  AC VDB(VO) PHASE(VO)
.PRINT  AC VDB(VD) PHASE(VD)
.PRINT  AC VDB(VIO) PHASE(VIO)
.PRINT  AC VDB(VGVG) PHASE(VGVG)
.PRINT  AC VDB(VGVD) PHASE(VGVD)
.PRINT  AC VDB(VIO2) PHASE(VIO2)
.PRINT  AC VDB(VI) PHASE(VI)
.PRINT  TRAN VO
.PRINT  TRAN VD
.PRINT  TRAN VIO
.PRINT  TRAN VGVG
.PRINT  TRAN VGVD
.PRINT  TRAN VIO2
.PRINT  TRAN VI
AGVG 1 5 LAPLACEA1
.MODEL LAPLACEA1 S_XFER( IN_OFFSET=0 GAIN=1 NUM_COEFF=[0.5]
+ DEN_COEFF=[7.8125E-9 2.5E-5 1] DENORM_FREQ=1)
AGVD 11 7 LAPLACEA2
.MODEL LAPLACEA2 S_XFER( IN_OFFSET=0 GAIN=1 NUM_COEFF=[10]
+ DEN_COEFF=[7.8125E-9 2.5E-5 1] DENORM_FREQ=1)
AZOUT 6 4 LAPLACEA3
.MODEL LAPLACEA3 S_XFER( IN_OFFSET=0 GAIN=1
+ NUM_COEFF=[125E-6 0] DEN_COEFF=[7.8125E-9 2.5E-5 1]
+ DENORM_FREQ=1)
VIO 6 0 DC=0 AC=0 PULSE 0 1 8M
VI 1 0 AC=0 PULSE 0 10 50U
X1 4 5 7 3 SUM3#0 
*{ K1=-1 K2=1 K3=1 }
.SUBCKT SUM3#0 1 2 3 4 
* 3 PORT SUMMER K1=GAIN1 K2=GAIN2 K3=GAIN3
B1 4 0 V = -1.0*V(1) + 1.0*V(2) + 1.0*V(3)
.ENDS
X2 14 2 8 SUM2#0 
*{ K1=-1 K2=1 }
.SUBCKT SUM2#0 1 2 3 
B1 3 0 V = -1.0*V(1) + 1.0*V(2)
.ENDS
XVM 9 11 GAIN#0 
*{ K=0.2 }
.SUBCKT GAIN#0 1 2
E1 2 0 1 0 200.0M
.ENDS
.SUBCKT GAIN#1 1 2
E1 2 0 1 0 500.0M
.ENDS
VREF 2 0 DC=2.5 AC=0
AGC 8 9 LAPLACEA6
.MODEL LAPLACEA6 S_XFER( IN_OFFSET=0 GAIN=1
+ NUM_COEFF=[0.03E-6 0.3427E-3 1] DEN_COEFF=[1.87E-15
+ 9.065E-10 0.17E-3 0] DENORM_FREQ=1)
XH 3 14 GAIN#1 
*{ K=0.5 }
.END
